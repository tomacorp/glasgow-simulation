* Translated from netlist ltspice/LM3880.cir
* /Users/toma/Documents/jitx/glasgow-simulation/model_lib/models/LM3880/ltspice/LM3880.asc
V1 VCC 0 PWL(0 0 100u 0 500u 5)
R2 EN 0 10K
V2 EN 0 PWL(0 0 100u 0 500u 1.15 1.5m 1.35 2m 5 3m 5 3.001m 0 10m 0 10.001m 3 160m 3 160.001m 0 240m 0 240.001m 3)
.tran 1u 320m
XLM3880 VCC 0 EN VCMPA VCMPB VCMPC LM3880
.subckt LM3880 VCC GND EN FLAG3 FLAG2 FLAG1
M1 VNI EN VSDP VSDP MDIFF
M2 VNP VZREF VSDP VSDP MDIFF
D1 GND VZREF DZREF
M3 VNI VNI VCC VCC MPMIR
M4 VNP VNP VCC VCC MPMIR
M5 ENA VNI VCC VCC MPGAIN
M6 ENB VNP VCC VCC MPGAIN
M7 VSDP GND GND GND MDISRC
M8 ENA VSG VSG VSG MDISRC
M9 ENB VSG VSG VSG MDISRC
M10 VCC VZREF VZREF VZREF MDISRC
R1 VCC EN 24.3K
M11 VSG GND GND GND MDIGAIN
M12 VCMP ENB VCC VCC MOSLOGP
M13 VCMP ENB GND GND MOSLOGN
M14 VCC EN EN EN MPPU
C1 EN GND 7pF
C2 VZREF GND 4pF
C3 ENB GND 1.3pF
C4 VNP GND 2.5pF
C5 VNI GND 2.5pF
C6 ENA GND 1.3pF
M15 VCMP GND VRGO VRGO MVREG
C7 VCMP GND 7pF
C8 VRGO GND 7pF
C9 VRAMP N003 5nF
D2 VRGI VRAMP DRAMP
M16 VDRMP VCMP VCMP VCMP MIRAMP
M17 VRGO VRGI VRGI VRGI MIRAMP
D3 VRAMP VDRMP DRAMP
C10 VDRMP VCMP 7pF
C11 VRGI VRGO 7pF
M18 VNIA VRAMP VSDPA VSDPA MDIFF
M19 VNPA VZREFA VSDPA VSDPA MDIFF
D4 GND VZREFA DZREFA
M20 VNIA VNIA VCC VCC MPMIR
M21 VNPA VNPA VCC VCC MPMIR
M22 ENAA VNPA VCC VCC MPGAIN
M23 ENBA VNIA VCC VCC MPGAIN
M24 VSDPA GND GND GND MDISRC
M25 ENAA VSGA VSGA VSGA MDISRC
M26 ENBA VSGA VSGA VSGA MDISRC
M27 VCC VZREFA VZREFA VZREFA MDISRC
M28 VSGA GND GND GND MDIGAIN
M29 FLAG3 ENAA VCC VCC MOSFLAGP
M30 FLAG3 ENAA GND GND MOSFLAGN
C13 VZREFA GND 4pF
C14 ENAA GND 1.3pF
C15 VNIA GND 2.5pF
C16 VNPA GND 2.5pF
C17 ENBA GND 1.3pF
C18 FLAG3 GND 7pF
M31 VNIB VRAMP VSDPB VSDPB MDIFF
M32 VNPB VZREFB VSDPB VSDPB MDIFF
D5 GND VZREFB DZREFB
M33 VNIB VNIB VCC VCC MPMIR
M34 VNPB VNPB VCC VCC MPMIR
M35 ENBB VNPB VCC VCC MPGAIN
M36 ENAB VNIB VCC VCC MPGAIN
M37 VSDPB GND GND GND MDISRC
M38 ENBB VSGB VSGB VSGB MDISRC
M39 ENAB VSGB VSGB VSGB MDISRC
M40 VCC VZREFB VZREFB VZREFB MDISRC
M41 VSGB GND GND GND MDIGAIN
M42 FLAG2 ENBB VCC VCC MOSFLAGP
M43 FLAG2 ENBB GND GND MOSFLAGN
C12 VZREFB GND 4pF
C19 ENBB GND 1.3pF
C20 VNIB GND 2.5pF
C21 VNPB GND 2.5pF
C22 ENAB GND 1.3pF
C23 FLAG2 GND 7pF
M44 VNIC VRAMP VSDPC VSDPC MDIFF
M45 VNPC VZREFC VSDPC VSDPC MDIFF
D6 GND VZREFC DZREFC
M46 VNIC VNIC VCC VCC MPMIR
M47 VNPC VNPC VCC VCC MPMIR
M48 ENAC VNPC VCC VCC MPGAIN
M49 N001 VNIC VCC VCC MPGAIN
M50 VSDPC GND GND GND MDISRC
M51 ENAC VSGC VSGC VSGC MDISRC
M52 N001 VSGC VSGC VSGC MDISRC
M53 VCC VZREFC VZREFC VZREFC MDISRC
M54 VSGC GND GND GND MDIGAIN
M55 FLAG1 ENAC VCC VCC MOSFLAGP
M56 FLAG1 ENAC GND GND MOSFLAGN
C24 VZREFC GND 4pF
C25 ENAC GND 1.3pF
C26 VNIC GND 2.5pF
C27 VNPC GND 2.5pF
C28 N001 GND 1.3pF
C29 FLAG1 GND 7pF
D7 GND EN DESD
D8 EN VCC DESD
D9 N003 VRAMP DZRAMP
M57 GND GND N003 N003 MPVN
C30 N003 GND 200pF
M59 VCC N003 N003 N003 MDISRC
.model MDIFF NMOS LEVEL=1 RD=10 RS=10 VTO=-0.35 KP=100u
.model MDISRC NMOS LEVEL=1 RD=10 RS=10 VTO=-0.35 KP=65.3u
.model MPMIR PMOS LEVEL=1 RD=10 RS=10 VTO=.35 KP=40u
.model MPGAIN PMOS LEVEL=1 RD=10 RS=10 VTO=0.15 KP=110u
.model MDIGAIN NMOS LEVEL=1 RD=10 RS=10 VTO=-0.35 KP=200u
.model MPPU NMOS LEVEL=1 RD=10 RS=10 VTO=-0.8 KP=21.875u
.model MOSLOGN NMOS LEVEL=1 RD=10 RS=10 VTO=0.8 KP=100u
.model MOSLOGP PMOS LEVEL=1 RD=10 RS=10 VTO=-0.3 KP=20u
.model MOSFLAGN NMOS LEVEL=1 RD=1 RS=1 VTO=0.8 KP=2.2m
.model MOSFLAGP PMOS LEVEL=1 RD=1 RS=1 VTO=-0.3 KP=440u
.model DZREF D RS=0.1 N=1 BV=1.25 IBV=4u
.model DZREFA D RS=0.1 N=1 BV=1.4 IBV=4u
.model DZREFB D RS=0.1 N=1 BV=1.1 IBV=4u
.model DZREFC D RS=0.1 N=1 BV=0.8 IBV=4u
.model DZRAMP D RS=0.1 N=1 BV=1.1 IBV=4u
.model DESD D RS=0.1 N=1 IS=1e-8
.model MVREG NMOS LEVEL=1 RD=10 RS=10 VTO=-2.2 KP=100u
.model MPVN PMOS LEVEL=1 RD=10 RS=10 VTO=-0.5 KP=10m
.model MIRAMP NMOS LEVEL=1 RD=10 RS=10 VTO=-0.5 KP=0.8u
.model DRAMP D RS=1000 N=1 IS=1e-12
.model QRAMP NPN BF=50 RE=1 RC=1 RB=10 CJE=10P
.ends
.end